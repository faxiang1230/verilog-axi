/*

Copyright (c) 2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * AXI4 RAM
 */
module axi_ram #
(
    // Width of data bus in bits
    parameter DATA_WIDTH = 32,
    // Width of address bus in bits
    parameter ADDR_WIDTH = 16,
    // Width of wstrb (width of data bus in words)
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    // Width of ID signal
    parameter ID_WIDTH = 8,
    // Extra pipeline register on output
    parameter PIPELINE_OUTPUT = 0,
    // Extra init file
    parameter INIT_FILE = ""
)
(
    input  wire                   clk,
    input  wire                   rst,

    input  wire [ID_WIDTH-1:0]    s_axi_awid,
    input  wire [ADDR_WIDTH-1:0]  s_axi_awaddr,
    input  wire [7:0]             s_axi_awlen,
    input  wire [2:0]             s_axi_awsize,
    input  wire [1:0]             s_axi_awburst,
    input  wire                   s_axi_awlock,
    input  wire [3:0]             s_axi_awcache,
    input  wire [2:0]             s_axi_awprot,
    input  wire                   s_axi_awvalid,
    output wire                   s_axi_awready,
    input  wire [DATA_WIDTH-1:0]  s_axi_wdata,
    input  wire [STRB_WIDTH-1:0]  s_axi_wstrb,
    input  wire                   s_axi_wlast,
    input  wire                   s_axi_wvalid,
    output wire                   s_axi_wready,
    output wire [ID_WIDTH-1:0]    s_axi_bid,
    output wire [1:0]             s_axi_bresp,
    output wire                   s_axi_bvalid,
    input  wire                   s_axi_bready,
    input  wire [ID_WIDTH-1:0]    s_axi_arid,
    input  wire [ADDR_WIDTH-1:0]  s_axi_araddr,
    input  wire [7:0]             s_axi_arlen,
    input  wire [2:0]             s_axi_arsize,
    input  wire [1:0]             s_axi_arburst,
    input  wire                   s_axi_arlock,
    input  wire [3:0]             s_axi_arcache,
    input  wire [2:0]             s_axi_arprot,
    input  wire                   s_axi_arvalid,
    output wire                   s_axi_arready,
    output wire [ID_WIDTH-1:0]    s_axi_rid,
    output wire [DATA_WIDTH-1:0]  s_axi_rdata,
    output wire [1:0]             s_axi_rresp,
    output wire                   s_axi_rlast,
    output wire                   s_axi_rvalid,
    input  wire                   s_axi_rready
);

parameter VALID_ADDR_WIDTH = ADDR_WIDTH - $clog2(STRB_WIDTH);
parameter WORD_WIDTH = STRB_WIDTH;
parameter WORD_SIZE = DATA_WIDTH/WORD_WIDTH;
localparam BUS_ADDR_WIDTH = $clog2(STRB_WIDTH);

// bus width assertions
initial begin
    if (WORD_SIZE * STRB_WIDTH != DATA_WIDTH) begin
        $error("Error: AXI data width not evenly divisble (instance %m)");
        $finish;
    end

    if (2**$clog2(WORD_WIDTH) != WORD_WIDTH) begin
        $error("Error: AXI word width must be even power of two (instance %m)");
        $finish;
    end
end

localparam [0:0]
    READ_STATE_IDLE = 1'd0,
    READ_STATE_BURST = 1'd1;

reg [0:0] read_state_reg = READ_STATE_IDLE, read_state_next;

localparam [1:0]
    WRITE_STATE_IDLE = 2'd0,
    WRITE_STATE_BURST = 2'd1,
    WRITE_STATE_RESP = 2'd2;

localparam [1:0]
	BURST_FIX  = 2'b00,
	BURST_INCR = 2'b01,
	BURST_WRAP = 2'b10;

reg [1:0] write_state_reg = WRITE_STATE_IDLE, write_state_next;

reg mem_wr_en;
reg mem_rd_en;

reg [ID_WIDTH-1:0] read_id_reg = {ID_WIDTH{1'b0}}, read_id_next;
reg [ADDR_WIDTH-1:0] read_addr_reg = {ADDR_WIDTH{1'b0}}, read_addr_next;
reg [7:0] read_count_reg = 8'd0, read_count_next;
reg [2:0] read_size_reg = 3'd0, read_size_next;
reg [1:0] read_burst_reg = 2'd0, read_burst_next;

reg [ADDR_WIDTH-1:12] read_wrap_high_addr_reg = {(ADDR_WIDTH-12){1'b0}}, read_wrap_high_addr_next;
reg [11:0] read_wrap_low_boundary_reg, read_wrap_low_boundary_next;
reg [11:0] read_wrap_high_boundary_reg, read_wrap_high_boundary_next;

reg [BUS_ADDR_WIDTH-1:0] read_wrap_low_addr_reg, read_wrap_low_addr_next;
reg [BUS_ADDR_WIDTH-1:0] read_wrap_low_align_addr_reg, read_wrap_low_align_addr_next;
reg [BUS_ADDR_WIDTH-1:0] read_wrap_low_addr_next_r1;

reg [11:BUS_ADDR_WIDTH] read_wrap_mid_addr_reg, read_wrap_mid_addr_next;
reg [11:BUS_ADDR_WIDTH] read_wrap_mid_addr_next_r1;
reg [11:0] read_wrap_mid_low_addr_next_r1;
reg read_wrap_low_addr_overflow, read_wrap_mid_addr_overflow;

reg [ID_WIDTH-1:0] write_id_reg = {ID_WIDTH{1'b0}}, write_id_next;
reg [ADDR_WIDTH-1:0] write_addr_reg = {ADDR_WIDTH{1'b0}}, write_addr_next;
reg [7:0] write_count_reg = 8'd0, write_count_next;
reg [2:0] write_size_reg = 3'd0, write_size_next;
reg [1:0] write_burst_reg = 2'd0, write_burst_next;

reg [ADDR_WIDTH-1:12] write_wrap_high_addr_reg = {(ADDR_WIDTH-12){1'b0}}, write_wrap_high_addr_next;
reg [11:0] write_wrap_low_boundary_reg, write_wrap_low_boundary_next;
reg [11:0] write_wrap_high_boundary_reg, write_wrap_high_boundary_next;

reg [BUS_ADDR_WIDTH-1:0] write_wrap_low_addr_reg, write_wrap_low_addr_next;
reg [BUS_ADDR_WIDTH-1:0] write_wrap_low_align_addr_reg, write_wrap_low_align_addr_next;
reg [BUS_ADDR_WIDTH-1:0] write_wrap_low_addr_next_r1;

reg [11:BUS_ADDR_WIDTH] write_wrap_mid_addr_reg, write_wrap_mid_addr_next;
reg [11:BUS_ADDR_WIDTH] write_wrap_mid_addr_next_r1;
reg [11:0] write_wrap_mid_low_addr_next_r1;
reg write_wrap_low_addr_overflow, write_wrap_mid_addr_overflow;

reg s_axi_awready_reg = 1'b0, s_axi_awready_next;
reg s_axi_wready_reg = 1'b0, s_axi_wready_next;
reg [ID_WIDTH-1:0] s_axi_bid_reg = {ID_WIDTH{1'b0}}, s_axi_bid_next;
reg s_axi_bvalid_reg = 1'b0, s_axi_bvalid_next;
reg s_axi_arready_reg = 1'b0, s_axi_arready_next;
reg [ID_WIDTH-1:0] s_axi_rid_reg = {ID_WIDTH{1'b0}}, s_axi_rid_next;
reg [DATA_WIDTH-1:0] s_axi_rdata_reg = {DATA_WIDTH{1'b0}}, s_axi_rdata_next;
reg s_axi_rlast_reg = 1'b0, s_axi_rlast_next;
reg s_axi_rvalid_reg = 1'b0, s_axi_rvalid_next;
reg [ID_WIDTH-1:0] s_axi_rid_pipe_reg = {ID_WIDTH{1'b0}};
reg [DATA_WIDTH-1:0] s_axi_rdata_pipe_reg = {DATA_WIDTH{1'b0}};
reg s_axi_rlast_pipe_reg = 1'b0;
reg s_axi_rvalid_pipe_reg = 1'b0;

// (* RAM_STYLE="BLOCK" *)
reg [DATA_WIDTH-1:0] mem[(2**VALID_ADDR_WIDTH)-1:0];

wire [VALID_ADDR_WIDTH-1:0] s_axi_awaddr_valid = s_axi_awaddr >> (ADDR_WIDTH - VALID_ADDR_WIDTH);
wire [VALID_ADDR_WIDTH-1:0] s_axi_araddr_valid = s_axi_araddr >> (ADDR_WIDTH - VALID_ADDR_WIDTH);
wire [VALID_ADDR_WIDTH-1:0] read_addr_valid = read_addr_reg >> (ADDR_WIDTH - VALID_ADDR_WIDTH);
wire [VALID_ADDR_WIDTH-1:0] write_addr_valid = write_addr_reg >> (ADDR_WIDTH - VALID_ADDR_WIDTH);

assign s_axi_awready = s_axi_awready_reg;
assign s_axi_wready = s_axi_wready_reg;
assign s_axi_bid = s_axi_bid_reg;
assign s_axi_bresp = 2'b00;
assign s_axi_bvalid = s_axi_bvalid_reg;
assign s_axi_arready = s_axi_arready_reg;
assign s_axi_rid = PIPELINE_OUTPUT ? s_axi_rid_pipe_reg : s_axi_rid_reg;
assign s_axi_rdata = PIPELINE_OUTPUT ? s_axi_rdata_pipe_reg : s_axi_rdata_reg;
assign s_axi_rresp = 2'b00;
assign s_axi_rlast = PIPELINE_OUTPUT ? s_axi_rlast_pipe_reg : s_axi_rlast_reg;
assign s_axi_rvalid = PIPELINE_OUTPUT ? s_axi_rvalid_pipe_reg : s_axi_rvalid_reg;

integer i, j;

initial begin
    // two nested loops for smaller number of iterations per loop
    // workaround for synthesizer complaints about large loop counts
    for (i = 0; i < 2**VALID_ADDR_WIDTH; i = i + 2**(VALID_ADDR_WIDTH/2)) begin
        for (j = i; j < i + 2**(VALID_ADDR_WIDTH/2); j = j + 1) begin
            mem[j] = 0;
        end
    end

    if (INIT_FILE != "") begin
       $readmemh(INIT_FILE, mem);
    end

end

always @* begin
    write_state_next = WRITE_STATE_IDLE;

    mem_wr_en = 1'b0;

    write_id_next = write_id_reg;
    write_addr_next = write_addr_reg;
    write_count_next = write_count_reg;
    write_size_next = write_size_reg;
    write_burst_next = write_burst_reg;

    s_axi_awready_next = 1'b0;
    s_axi_wready_next = 1'b0;
    s_axi_bid_next = s_axi_bid_reg;
    s_axi_bvalid_next = s_axi_bvalid_reg && !s_axi_bready;

    write_wrap_high_addr_next = write_wrap_high_addr_reg;
    write_wrap_mid_addr_next = write_wrap_mid_addr_reg;
    write_wrap_low_addr_next = write_wrap_low_addr_reg;
    write_wrap_low_align_addr_next = write_wrap_low_align_addr_reg;

    write_wrap_low_boundary_next = write_wrap_low_boundary_reg;
    write_wrap_high_boundary_next = write_wrap_high_boundary_reg;
    write_wrap_low_addr_overflow = 1'b0;
    write_wrap_mid_addr_overflow = 1'b0;

    case (write_state_reg)
        WRITE_STATE_IDLE: begin
            s_axi_awready_next = 1'b1;

            if (s_axi_awready && s_axi_awvalid) begin
                write_id_next = s_axi_awid;
                write_addr_next = s_axi_awaddr;
                write_count_next = s_axi_awlen;
                write_size_next = s_axi_awsize < $clog2(STRB_WIDTH) ? s_axi_awsize : $clog2(STRB_WIDTH);
                write_burst_next = s_axi_awburst;

                write_wrap_high_addr_next = s_axi_awaddr[ADDR_WIDTH-1:12];
                write_wrap_mid_addr_next = s_axi_awaddr[11:BUS_ADDR_WIDTH];
                write_wrap_low_addr_next = s_axi_awaddr[BUS_ADDR_WIDTH-1:0];

                write_wrap_low_align_addr_next = s_axi_awaddr[BUS_ADDR_WIDTH-1:0] &
                    ({BUS_ADDR_WIDTH{1'b1}} & ~((1 << write_size_next) - 1));
                write_wrap_low_boundary_next = s_axi_awaddr[11:0] & ~(((s_axi_awlen[3:0] + 1) << write_size_next) - 1);
                write_wrap_high_boundary_next = write_wrap_low_boundary_next + ((s_axi_awlen[3:0] + 1) << write_size_next);

                s_axi_awready_next = 1'b0;
                s_axi_wready_next = 1'b1;
                write_state_next = WRITE_STATE_BURST;
            end else begin
                write_state_next = WRITE_STATE_IDLE;
            end
        end
        WRITE_STATE_BURST: begin
            s_axi_wready_next = 1'b1;

            if (s_axi_wready && s_axi_wvalid) begin
                mem_wr_en = 1'b1;
                if (write_burst_reg == BURST_INCR) begin
                    write_addr_next = write_addr_reg + (1 << write_size_reg);
				end else if (write_burst_reg == BURST_WRAP) begin
                    {write_wrap_low_addr_overflow, write_wrap_low_addr_next_r1} = write_wrap_low_align_addr_reg + (1 << write_size_reg);
                    {write_wrap_mid_addr_overflow, write_wrap_mid_addr_next_r1} = write_wrap_mid_addr_reg + 1;

                    write_wrap_mid_low_addr_next_r1 = write_wrap_low_addr_overflow ?
                        {write_wrap_mid_addr_next_r1, write_wrap_low_addr_next_r1}:
                        {write_wrap_mid_addr_reg, write_wrap_low_addr_next_r1};

                    write_addr_next = (write_wrap_mid_low_addr_next_r1 == write_wrap_high_boundary_reg) ?
                        {write_wrap_high_addr_reg, write_wrap_low_boundary_reg} :
                        {write_wrap_high_addr_reg, write_wrap_mid_low_addr_next_r1};

                    write_wrap_low_align_addr_next = write_addr_next[BUS_ADDR_WIDTH-1:0];
                end
                write_count_next = write_count_reg - 1;
                if (write_count_reg > 0) begin
                    write_state_next = WRITE_STATE_BURST;
                end else begin
                    s_axi_wready_next = 1'b0;
                    if (s_axi_bready || !s_axi_bvalid) begin
                        s_axi_bid_next = write_id_reg;
                        s_axi_bvalid_next = 1'b1;
                        s_axi_awready_next = 1'b1;
                        write_state_next = WRITE_STATE_IDLE;
                    end else begin
                        write_state_next = WRITE_STATE_RESP;
                    end
                end
            end else begin
                write_state_next = WRITE_STATE_BURST;
            end
        end
        WRITE_STATE_RESP: begin
            if (s_axi_bready || !s_axi_bvalid) begin
                s_axi_bid_next = write_id_reg;
                s_axi_bvalid_next = 1'b1;
                s_axi_awready_next = 1'b1;
                write_state_next = WRITE_STATE_IDLE;
            end else begin
                write_state_next = WRITE_STATE_RESP;
            end
        end
    endcase
end

always @(posedge clk) begin
    write_state_reg <= write_state_next;

    write_id_reg <= write_id_next;
    write_addr_reg <= write_addr_next;
    write_count_reg <= write_count_next;
    write_size_reg <= write_size_next;
    write_burst_reg <= write_burst_next;

    s_axi_awready_reg <= s_axi_awready_next;
    s_axi_wready_reg <= s_axi_wready_next;
    s_axi_bid_reg <= s_axi_bid_next;
    s_axi_bvalid_reg <= s_axi_bvalid_next;

    write_wrap_high_addr_reg <= write_wrap_high_addr_next;
    write_wrap_mid_addr_reg <= write_addr_next[11:BUS_ADDR_WIDTH];
    write_wrap_low_addr_reg <= write_addr_next[BUS_ADDR_WIDTH-1:0];
    write_wrap_low_align_addr_reg <= write_wrap_low_align_addr_next;
    write_wrap_low_boundary_reg <= write_wrap_low_boundary_next;
    write_wrap_high_boundary_reg <= write_wrap_high_boundary_next;

    for (i = 0; i < WORD_WIDTH; i = i + 1) begin
        if (mem_wr_en & s_axi_wstrb[i]) begin
            mem[write_addr_valid][WORD_SIZE*i +: WORD_SIZE] <= s_axi_wdata[WORD_SIZE*i +: WORD_SIZE];
        end
    end

    if (rst) begin
        write_state_reg <= WRITE_STATE_IDLE;

        s_axi_awready_reg <= 1'b0;
        s_axi_wready_reg <= 1'b0;
        s_axi_bvalid_reg <= 1'b0;
    end
end

always @* begin
    read_state_next = READ_STATE_IDLE;

    mem_rd_en = 1'b0;

    s_axi_rid_next = s_axi_rid_reg;
    s_axi_rlast_next = s_axi_rlast_reg;
    s_axi_rvalid_next = s_axi_rvalid_reg && !(s_axi_rready || (PIPELINE_OUTPUT && !s_axi_rvalid_pipe_reg));

    read_id_next = read_id_reg;
    read_addr_next = read_addr_reg;
    read_count_next = read_count_reg;
    read_size_next = read_size_reg;
    read_burst_next = read_burst_reg;

    read_wrap_high_addr_next = read_wrap_high_addr_reg;
    read_wrap_mid_addr_next = read_wrap_mid_addr_reg;
    read_wrap_low_addr_next = read_wrap_low_addr_reg;
    read_wrap_low_align_addr_next = read_wrap_low_align_addr_reg;

    read_wrap_low_boundary_next = read_wrap_low_boundary_reg;
    read_wrap_high_boundary_next = read_wrap_high_boundary_reg;
    read_wrap_low_addr_overflow = 1'b0;
    read_wrap_mid_addr_overflow = 1'b0;

    s_axi_arready_next = 1'b0;

    case (read_state_reg)
        READ_STATE_IDLE: begin
            s_axi_arready_next = 1'b1;
            s_axi_rlast_next = 1'b0;

            if (s_axi_arready && s_axi_arvalid) begin
                read_id_next = s_axi_arid;
                read_addr_next = s_axi_araddr;
                read_count_next = s_axi_arlen;
                read_size_next = s_axi_arsize < $clog2(STRB_WIDTH) ? s_axi_arsize : $clog2(STRB_WIDTH);
                read_burst_next = s_axi_arburst;

                read_wrap_high_addr_next = s_axi_araddr[ADDR_WIDTH-1:12];
                read_wrap_mid_addr_next = s_axi_araddr[11:BUS_ADDR_WIDTH];
                read_wrap_low_addr_next = s_axi_araddr[BUS_ADDR_WIDTH-1:0];

                read_wrap_low_align_addr_next = s_axi_araddr[BUS_ADDR_WIDTH-1:0] &
                    ({BUS_ADDR_WIDTH{1'b1}} & ~((1 << read_size_next) - 1));
                read_wrap_low_boundary_next = s_axi_araddr[11:0] & ~(((s_axi_arlen[3:0] + 1) << read_size_next) - 1);
                read_wrap_high_boundary_next = read_wrap_low_boundary_next + ((s_axi_arlen[3:0] + 1) << read_size_next);

                s_axi_arready_next = 1'b0;
                read_state_next = READ_STATE_BURST;
            end else begin
                read_state_next = READ_STATE_IDLE;
            end
        end
        READ_STATE_BURST: begin
            if (s_axi_rready || (PIPELINE_OUTPUT && !s_axi_rvalid_pipe_reg) || !s_axi_rvalid_reg) begin
                mem_rd_en = 1'b1;
                s_axi_rvalid_next = 1'b1;
                s_axi_rid_next = read_id_reg;
                s_axi_rlast_next = read_count_reg == 0;
                if (read_burst_reg == BURST_INCR) begin
                    read_addr_next = read_addr_reg + (1 << read_size_reg);
                end else if (read_burst_reg == BURST_WRAP) begin
                    {read_wrap_low_addr_overflow, read_wrap_low_addr_next_r1} = read_wrap_low_align_addr_reg + (1 << read_size_reg);
                    {read_wrap_mid_addr_overflow, read_wrap_mid_addr_next_r1} = read_wrap_mid_addr_reg + 1;

                    read_wrap_mid_low_addr_next_r1 = read_wrap_low_addr_overflow ?
                        {read_wrap_mid_addr_next_r1, read_wrap_low_addr_next_r1}:
                        {read_wrap_mid_addr_reg, read_wrap_low_addr_next_r1};

                    read_addr_next = (read_wrap_mid_low_addr_next_r1 == read_wrap_high_boundary_reg) ?
                        {read_wrap_high_addr_reg, read_wrap_low_boundary_reg} :
                        {read_wrap_high_addr_reg, read_wrap_mid_low_addr_next_r1};

                    read_wrap_low_align_addr_next = read_addr_next[BUS_ADDR_WIDTH-1:0];
                end
                read_count_next = read_count_reg - 1;
                if (read_count_reg > 0) begin
                    read_state_next = READ_STATE_BURST;
                end else begin
                    s_axi_arready_next = 1'b1;
                    read_state_next = READ_STATE_IDLE;
                end
            end else begin
                read_state_next = READ_STATE_BURST;
            end
        end
    endcase
end

always @(posedge clk) begin
    read_state_reg <= read_state_next;

    read_id_reg <= read_id_next;
    read_addr_reg <= read_addr_next;
    read_count_reg <= read_count_next;
    read_size_reg <= read_size_next;
    read_burst_reg <= read_burst_next;

    s_axi_arready_reg <= s_axi_arready_next;
    s_axi_rid_reg <= s_axi_rid_next;
    s_axi_rlast_reg <= s_axi_rlast_next;
    s_axi_rvalid_reg <= s_axi_rvalid_next;

    read_wrap_high_addr_reg <= read_wrap_high_addr_next;
    read_wrap_mid_addr_reg <= read_addr_next[11:BUS_ADDR_WIDTH];
    read_wrap_low_addr_reg <= read_addr_next[BUS_ADDR_WIDTH-1:0];
    read_wrap_low_align_addr_reg <= read_wrap_low_align_addr_next;
    read_wrap_low_boundary_reg <= read_wrap_low_boundary_next;
    read_wrap_high_boundary_reg <= read_wrap_high_boundary_next;

    if (mem_rd_en) begin
        s_axi_rdata_reg <= mem[read_addr_valid];
    end

    if (!s_axi_rvalid_pipe_reg || s_axi_rready) begin
        s_axi_rid_pipe_reg <= s_axi_rid_reg;
        s_axi_rdata_pipe_reg <= s_axi_rdata_reg;
        s_axi_rlast_pipe_reg <= s_axi_rlast_reg;
        s_axi_rvalid_pipe_reg <= s_axi_rvalid_reg;
    end

    if (rst) begin
        read_state_reg <= READ_STATE_IDLE;

        s_axi_arready_reg <= 1'b0;
        s_axi_rvalid_reg <= 1'b0;
        s_axi_rvalid_pipe_reg <= 1'b0;
    end
end

endmodule

`resetall
